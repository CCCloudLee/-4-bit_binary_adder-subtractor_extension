//???_E94084016
//implement 4-bit adder
module four_bit_full_adder (sum, Cout, a, b, Cin);
  input [3:0] a;
  input [3:0] b;
  input Cin; //carry in
  output [3:0] sum;
  output Cout; //carry out
  wire [3:0] c;

  one_bit_full_adder fa1(sum[0], c[1], a[0],b[0], Cin ) ;
  one_bit_full_adder fa2(sum[1], c[2], a[1],b[1], c[1] ) ;
  one_bit_full_adder fa3(sum[2], c[3], a[2],b[2], c[2] ) ;
  one_bit_full_adder fa4(sum[3], Cout, a[3],b[3], c[3] ) ;

endmodule